module not_16(
  input wire [15:0] in,
  output wire [15:0] out
);
  not_0 n0(in[0], out[0]);
  not_0 n1(in[1], out[1]);
  not_0 n2(in[2], out[2]);
  not_0 n3(in[3], out[3]);
  not_0 n4(in[4], out[4]);
  not_0 n5(in[5], out[5]);
  not_0 n6(in[6], out[6]);
  not_0 n7(in[7], out[7]);
  not_0 n8(in[8], out[8]);
  not_0 n9(in[9], out[9]);
  not_0 n10(in[10], out[10]);
  not_0 n11(in[11], out[11]);
  not_0 n12(in[12], out[12]);
  not_0 n13(in[13], out[13]);
  not_0 n14(in[14], out[14]);
  not_0 n15(in[15], out[15]);
endmodule
