module alu(
  input wire x[15:0],
  input wire y[15:0],
  input wire zx,
  input wire nx,
  input wire zy,
  input wire ny,
  input wire f,
  input wire no,
  output wire out[15:0],
  output wire zr,
  output wire ng
);
endmodule
