`include "testbench/assert.v"

module or_16_testbench;
  reg [15:0] a, b;
  wire [15:0] out;

  or_16 o16(a, b, out);

  initial begin
    a=16'b0000000000000000;
    b=16'b0000000000000000;
    #10;
    `assert(out, 16'b0000000000000000);

    a=16'b0000000000000000;
    b=16'b1111111111111111;
    #10;
    `assert(out, 16'b1111111111111111);

    a=16'b1111111111111111;
    b=16'b1111111111111111;
    #10;
    `assert(out, 16'b1111111111111111);

    a=16'b1010101010101010;
    b=16'b0101010101010101;
    #10;
    `assert(out, 16'b1111111111111111);

    a=16'b0011110011000011;
    b=16'b0000111111110000;
    #10;
    `assert(out, 16'b0011111111110011);

    a=16'b0001001000110100;
    b=16'b1001100001110110;
    #10;
    `assert(out, 16'b1001101001110110);
  end
endmodule
